module M_WB_register (
    input 
);
    
endmodule