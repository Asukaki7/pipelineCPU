module EX_Mul3BusBFW (
    //control port
    input [1:0] BusBFW,

    //input data
    input [31:0] busB_EX,
    input [31:0] Di,
    input [31:0] ALUout_M,
    

    output reg [31:0] BusBFW_out
);

always @(*) begin
    case (BusBFW)
        2'b00: begin
            BusBFW_out <= busB_EX;
        end 

        2'b01:begin
            BusBFW_out <= Di;
        end

        2'b10:begin
            BusBFW_out <= ALUout_M;
        end
        
        default:begin
            BusBFW_out <= 32'h0000_0000;
        end 
    endcase
end


endmodule