module ID(
    
);


endmodule